LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-----------------------------------------------------
ENTITY uProgramMemory IS
PORT(	uaddr	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
		UI		: 	OUT 	STD_LOGIC_VECTOR(28 DOWNTO 0));
END ENTITY uProgramMemory;
-----------------------------------------------------
ARCHITECTURE behavioral OF uProgramMemory IS
BEGIN
	
	MUI: PROCESS(uaddr)
	BEGIN
		CASE uaddr IS
	-- Complete the following values according to your particular implementation 
	-- Unused postions do not affect the operation of the ROM
			-- FETCH 							    
			WHEN "00000000" => UI <= "00000000100001000000010110101"; 
			WHEN "00000001" => UI <= "00000000000001000000010000000"; 
			WHEN "00000010" => UI <= "01100000000010000000010000000"; 
			WHEN "00000011" => UI <= "00000000000000110000010000000"; 
			WHEN "00000100" => UI <= "00000000000000010001011000000";
		
			-- INT
			WHEN "00000101" => UI <= "00000000000000101000010000000"; 
			WHEN "00000110" => UI <= "01100000100110000010010000000"; 
			WHEN "00000111" => UI <= "00010010000010000001111000000"; 

			--00001	 MOV ACC,A 
			WHEN "00001000" => UI <= "10000001111110000001111000000";
			WHEN "00001001" => UI <= "00000000000000000000000000000";
			WHEN "00001010" => UI <= "00000000000000000000000000000";
			WHEN "00001011" => UI <= "00000000000000000000000000000";
			WHEN "00001100" => UI <= "00000000000000000000000000000";
			WHEN "00001101" => UI <= "00000000000000000000000000000";
			WHEN "00001110" => UI <= "00000000000000000000000000000";
			WHEN "00001111" => UI <= "00000000000000000000000000000";

			--00010  MOV A,ACC
			WHEN "00010000" => UI <= "10000011101110000001111000000";
			WHEN "00010001" => UI <= "00000000000000000000000000000";
			WHEN "00010010" => UI <= "00000000000000000000000000000";
			WHEN "00010011" => UI <= "00000000000000000000000000000";
			WHEN "00010100" => UI <= "00000000000000000000000000000";
			WHEN "00010101" => UI <= "00000000000000000000000000000";
			WHEN "00010110" => UI <= "00000000000000000000000000000";
			WHEN "00010111" => UI <= "00000000000000000000000000000";

			--00011	 MOV ACC,CTE
			WHEN "00011000" => UI <= "00000000011101000000010000000";
			WHEN "00011001" => UI <= "01100000000010000000010000000";
			WHEN "00011010" => UI <= "00000000011100110000010000000";
			WHEN "00011011" => UI <= "00000000011110010001111000000";
			WHEN "00011100" => UI <= "00000000000000000000000000000";
			WHEN "00011101" => UI <= "00000000000000000000000000000";
			WHEN "00011110" => UI <= "00000000000000000000000000000";
			WHEN "00011111" => UI <= "00000000000000000000000000000";

			--00100  MOV ACC,[DPTR]
			WHEN "00100000" => UI <= "00000001011101000000010000000";
			WHEN "00100001" => UI <= "00000001011100000000010000000";
			WHEN "00100010" => UI <= "00000001011100110000010000000";
			WHEN "00100011" => UI <= "00000001011110010001111000000";
			WHEN "00100100" => UI <= "00000000000000000000000000000";
			WHEN "00100101" => UI <= "00000000000000000000000000000";
			WHEN "00100110" => UI <= "00000000000000000000000000000";
			WHEN "00100111" => UI <= "00000000000000000000000000000";

			--00101  MOV DPTR,ACC
			WHEN "00101000" => UI <= "10000011101010000001111000000";
			WHEN "00101001" => UI <= "00000000000000000000000000000";
			WHEN "00101010" => UI <= "00000000000000000000000000000";
			WHEN "00101011" => UI <= "00000000000000000000000000000";
			WHEN "00101100" => UI <= "00000000000000000000000000000";
			WHEN "00101101" => UI <= "00000000000000000000000000000";
			WHEN "00101110" => UI <= "00000000000000000000000000000";
			WHEN "00101111" => UI <= "00000000000000000000000000000";

			-- 00110 MOV [DPTR],ACC	
			WHEN "00110000" => UI <= "00000001011101000000010000000";
			WHEN "00110001" => UI <= "00000011111100100000010000000";
			WHEN "00110010" => UI <= "10000011111100000011111000000";
			WHEN "00110011" => UI <= "00000000000000000000000000000";
			WHEN "00110100" => UI <= "00000000000000000000000000000";
			WHEN "00110101" => UI <= "00000000000000000000000000000";
			WHEN "00110110" => UI <= "00000000000000000000000000000";
			WHEN "00110111" => UI <= "00000000000000000000000000000";

			-- 00111 INV ACC
			WHEN "00111000" => UI <= "10010011111110000001111000000";
			WHEN "00111001" => UI <= "00000000000000000000000000000";
			WHEN "00111010" => UI <= "00000000000000000000000000000";
			WHEN "00111011" => UI <= "00000000000000000000000000000";
			WHEN "00111100" => UI <= "00000000000000000000000000000";
			WHEN "00111101" => UI <= "00000000000000000000000000000";
			WHEN "00111110" => UI <= "00000000000000000000000000000";
			WHEN "00111111" => UI <= "00000000000000000000000000000";
			
			 -- 01000 AND ACC,A	 
			WHEN "01000000" => UI <= "10100001111110000001111000000";
			WHEN "01000001" => UI <= "00000000000000000000000000000";
			WHEN "01000010" => UI <= "00000000000000000000000000000";
			WHEN "01000011" => UI <= "00000000000000000000000000000";
			WHEN "01000100" => UI <= "00000000000000000000000000000";
			WHEN "01000101" => UI <= "00000000000000000000000000000";
			WHEN "01000110" => UI <= "00000000000000000000000000000";
			WHEN "01000111" => UI <= "00000000000000000000000000000";
			
			-- 01001 ADD ACC,A
			WHEN "01001000" => UI <= "11010001111110000001111000000";
			WHEN "01001001" => UI <= "00000000000000000000000000000";
			WHEN "01001010" => UI <= "00000000000000000000000000000";
			WHEN "01001011" => UI <= "00000000000000000000000000000";
			WHEN "01001100" => UI <= "00000000000000000000000000000";
			WHEN "01001101" => UI <= "00000000000000000000000000000";
			WHEN "01001110" => UI <= "00000000000000000000000000000";
			WHEN "01001111" => UI <= "00000000000000000000000000000";
			
			-- 01010 JMP DIR
			WHEN "01010000" => UI <= "00000000000001000000010001010";
			WHEN "01010001" => UI <= "01100000000010000001111000000";
			WHEN "01010010" => UI <= "00000000000000000000010000000";
			WHEN "01010011" => UI <= "00000000000000100000010000000";
			WHEN "01010100" => UI <= "00000000000010010001111000000";
			WHEN "01010101" => UI <= "00000000000000000000000000000";
			WHEN "01010110" => UI <= "00000000000000000000000000000";
			WHEN "01010111" => UI <= "00000000000000000000000000000";
			
			-- 01011 JZ DIR
			WHEN "01011000" => UI <= "00000000000001000000010010010";
			WHEN "01011001" => UI <= "01100000000010000001111000000";
			WHEN "01011010" => UI <= "00000000000000000000010000000";
			WHEN "01011011" => UI <= "00000000000000100000010000000";
			WHEN "01011100" => UI <= "00000000000010010001111000000";
			WHEN "01011101" => UI <= "00000000000000000000000000000";
			WHEN "01011110" => UI <= "00000000000000000000000000000";
			WHEN "01011111" => UI <= "00000000000000000000000000000";

			-- 01100 JN DIR
			WHEN "01100000" => UI <= "00000000000001000000010011010";
			WHEN "01100001" => UI <= "01100000000010000001111000000";
			WHEN "01100010" => UI <= "00000000000000000000010000000";
			WHEN "01100011" => UI <= "00000000000000100000010000000";
			WHEN "01100100" => UI <= "00000000000010010001111000000";
			WHEN "01100101" => UI <= "00000000000000000000000000000";
			WHEN "01100110" => UI <= "00000000000000000000000000000";
			WHEN "01100111" => UI <= "00000000000000000000000000000";
			
			-- 01101 JC DIR
			WHEN "01101000" => UI <= "00000000000001000000010100010";
			WHEN "01101001" => UI <= "01100000000010000001111000000";
			WHEN "01101010" => UI <= "00000000000000000000010000000";
			WHEN "01101011" => UI <= "00000000000000100000010000000";
			WHEN "01101100" => UI <= "00000000000010010001111000000";
			WHEN "01101101" => UI <= "00000000000000000000000000000";
			WHEN "01101110" => UI <= "00000000000000000000000000000";
			WHEN "01101111" => UI <= "00000000000000000000000000000";
			
			-- 01110  CALL DIR       
			WHEN "01110000" => UI <= "00000000100001000000010000000";
			WHEN "01110001" => UI <= "01100000000000100001111000000";
			WHEN "01110010" => UI <= "01100000100110000010010000000";
			WHEN "01110011" => UI <= "00000000000001000000010000000";
			WHEN "01110100" => UI <= "00000000000000000000010000000";
			WHEN "01110101" => UI <= "00000000000000100000010000000";
			WHEN "01110110" => UI <= "00000000000010010001111000000";
			WHEN "01110111" => UI <= "00000000000000000000000000000";
			
			
			-- 01111  RET
			WHEN "01111000" => UI <= "00000011110110000000010000000";
			WHEN "01111001" => UI <= "00000000111110000000010000000";
			WHEN "01111010" => UI <= "01010011000111000000010000000";
			WHEN "01111011" => UI <= "00000000000000000000010000000";
			WHEN "01111100" => UI <= "00000000000000100000010000000";
			WHEN "01111101" => UI <= "00000000000010010000010000000";
			WHEN "01111110" => UI <= "00000010111110000001111000000";
			WHEN "01111111" => UI <= "00000000000000000000000000000";

			-- 10000  OR ACC,A
			WHEN "10000000" => UI <= "10110001111110000001111000000";
			WHEN "10000001" => UI <= "00000000000000000000000000000";
			WHEN "10000010" => UI <= "00000000000000000000000000000";
			WHEN "10000011" => UI <= "00000000000000000000000000000";
			WHEN "10000100" => UI <= "00000000000000000000000000000";
			WHEN "10000101" => UI <= "00000000000000000000000000000";
			WHEN "10000110" => UI <= "00000000000000000000000000000";
			WHEN "10000111" => UI <= "00000000000000000000000000000";
			
			-- 10001  XOR ACC,A
			WHEN "10001000" => UI <= "11000001111110000001111000000";
			WHEN "10001001" => UI <= "00000000000000000000000000000";
			WHEN "10001010" => UI <= "00000000000000000000000000000";
			WHEN "10001011" => UI <= "00000000000000000000000000000";
			WHEN "10001100" => UI <= "00000000000000000000000000000";
			WHEN "10001101" => UI <= "00000000000000000000000000000";
			WHEN "10001110" => UI <= "00000000000000000000000000000";
			WHEN "10001111" => UI <= "00000000000000000000000000000";
			
			-- 10010  INC ACC
			WHEN "10010000" => UI <= "11100011111110000001111000000";
			WHEN "10010001" => UI <= "00000000000000000000000000000";
			WHEN "10010010" => UI <= "00000000000000000000000000000";
			WHEN "10010011" => UI <= "00000000000000000000000000000";
			WHEN "10010100" => UI <= "00000000000000000000000000000";
			WHEN "10010101" => UI <= "00000000000000000000000000000";
			WHEN "10010110" => UI <= "00000000000000000000000000000";
			WHEN "10010111" => UI <= "00000000000000000000000000000";
			
			-- 10011  NEG ACC
			WHEN "10011000" => UI <= "11110011111110000001111000000";
			WHEN "10011001" => UI <= "00000000000000000000000000000";
			WHEN "10011010" => UI <= "00000000000000000000000000000";
			WHEN "10011011" => UI <= "00000000000000000000000000000";
			WHEN "10011100" => UI <= "00000000000000000000000000000";
			WHEN "10011101" => UI <= "00000000000000000000000000000";
			WHEN "10011110" => UI <= "00000000000000000000000000000";
			WHEN "10011111" => UI <= "00000000000000000000000000000";
			
			-- 10100  SLL ACC
			WHEN "10100000" => UI <= "00001011111110000001111000000";
			WHEN "10100001" => UI <= "00000000000000000000000000000";
			WHEN "10100010" => UI <= "00000000000000000000000000000";
			WHEN "10100011" => UI <= "00000000000000000000000000000";
			WHEN "10100100" => UI <= "00000000000000000000000000000";
			WHEN "10100101" => UI <= "00000000000000000000000000000";
			WHEN "10100110" => UI <= "00000000000000000000000000000";
			WHEN "10100111" => UI <= "00000000000000000000000000000";
			
			-- 10101  SLR ACC
			WHEN "10101000" => UI <= "00000111111110000001111000000";
			WHEN "10101001" => UI <= "00000000000000000000000000000";
			WHEN "10101010" => UI <= "00000000000000000000000000000";
			WHEN "10101011" => UI <= "00000000000000000000000000000";
			WHEN "10101100" => UI <= "00000000000000000000000000000";
			WHEN "10101101" => UI <= "00000000000000000000000000000";
			WHEN "10101110" => UI <= "00000000000000000000000000000";
			WHEN "10101111" => UI <= "00000000000000000000000000000";
			
			-- 10110  HALT
			WHEN "10110000" => UI <= "00000000000000000000000000000";
			WHEN "10110001" => UI <= "00000000000000000000000000000";
			WHEN "10110010" => UI <= "00000000000000000000000000000";
			WHEN "10110011" => UI <= "00000000000000000000000000000";
			WHEN "10110100" => UI <= "00000000000000000000000000000";
			WHEN "10110101" => UI <= "00000000000000000000000000000";
			WHEN "10110110" => UI <= "00000000000000000000000000000";
			WHEN "10110111" => UI <= "00000000000000000000000000000";
			
								
			------------------------------------
			-- Unused cases:
			WHEN others => UI <= (others => 'X');
		END CASE;
	END PROCESS;
END ARCHITECTURE Behavioral;



